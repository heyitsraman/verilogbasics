//Tak_01 Hello World Example
module hello_world ();

//Display message in console on a new line with tab before
initial begin
    $display("\n\t Hello World! \n");
    $display("\n\t End of the task! \n");        //Added another text after first simulation
end
    
endmodule
